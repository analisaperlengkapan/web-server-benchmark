module main

import vweb
import json

struct App {
	vweb.Context
}

@['/hello']
pub fn (mut app App) hello() vweb.Result {
	app.set_content_type('application/json')
	response := json.encode({'message': 'Hello, world!'})
	return app.text(response)
}

fn main() {
	mut app := &App{}
	vweb.run(app, 8080)
}
